library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Package_CB_Configuration is

-- Declare constants

  	constant CBCrystalsCount : integer := 720;
	constant CBNeighboursCount : integer := 12;

	--upwards or downwards crystal
	constant CBCrystalsOrientation : STD_LOGIC_VECTOR(0 to CBCrystalsCount-1) := "101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010101100101011001010110010";
	--belongs the Crystal to one of the 10 pole crystals (category 3 and 4)?
   constant CBCrystalsIsPole : STD_LOGIC_VECTOR(0 to CBCrystalsCount-1) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
	-- only '1' for crystal 5/1/1 and 4/1/1 for rule 2.5.1
   constant CBCrystalsIsOnly2Pole : STD_LOGIC_VECTOR(0 to CBCrystalsCount-1) := "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	--belongs the Crystal to category 6 and 7?
   constant CBCrystalsIsCutEdge : STD_LOGIC_VECTOR(0 to CBCrystalsCount-1) := "101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100100001001101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100100001001101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100100001001101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100100001001101000001010000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000100100001001";
	type Type_CrystalNeighbours is array(0 to CBCrystalsCount-1, 1 to CBNeighboursCount) of integer;
	constant CBCrystalNeighbours : Type_CrystalNeighbours := ( 
(576, 144, 1, 577, 432, 288, 145, 3, 2, 576, 146, 579), 
(3, 2, 0, 146, 4, 5, 579, 576, 144, 6, 577, 145), 
(579, 1, 5, 580, 577, 0, 3, 6, 8, 576, 4, 624), 
(1, 146, 4, 2, 0, 145, 149, 48, 6, 144, 152, 5), 
(48, 6, 3, 152, 49, 7, 5, 1, 146, 50, 2, 149), 
(6, 8, 2, 4, 7, 9, 624, 579, 1, 11, 580, 3), 
(5, 4, 7, 8, 2, 3, 48, 50, 11, 1, 49, 9), 
(50, 11, 6, 49, 53, 12, 9, 5, 4, 56, 8, 48), 
(624, 5, 9, 625, 580, 2, 6, 11, 10, 579, 7, 627), 
(11, 10, 8, 7, 12, 13, 627, 624, 5, 14, 625, 6), 
(627, 9, 13, 628, 625, 8, 11, 14, 16, 624, 12, 672), 
(9, 7, 12, 10, 8, 6, 50, 56, 14, 5, 53, 13), 
(56, 14, 11, 53, 57, 15, 13, 9, 7, 58, 10, 50), 
(14, 16, 10, 12, 15, 17, 672, 627, 9, 19, 628, 11), 
(13, 12, 15, 16, 10, 11, 56, 58, 19, 9, 57, 17), 
(58, 19, 14, 57, 61, 20, 17, 13, 12, 64, 16, 56), 
(672, 13, 17, 673, 628, 10, 14, 19, 18, 627, 15, 675), 
(19, 18, 16, 15, 20, 21, 675, 672, 13, 22, 673, 14), 
(675, 17, 21, 676, 673, 16, 19, 22, 24, 672, 20, 24), 
(17, 15, 20, 18, 16, 14, 58, 64, 22, 13, 61, 21), 
(64, 22, 19, 61, 65, 23, 21, 17, 15, 66, 18, 58), 
(22, 24, 18, 20, 23, 25, 676, 675, 17, 27, 675, 19), 
(21, 20, 23, 24, 18, 19, 64, 66, 27, 17, 65, 25), 
(66, 27, 22, 65, 69, 28, 25, 21, 20, 72, 24, 64), 
(676, 21, 25, 678, 675, 18, 22, 27, 26, 18, 23, 679), 
(27, 26, 24, 23, 28, 29, 679, 676, 21, 30, 678, 22), 
(679, 25, 29, 683, 678, 24, 27, 30, 32, 676, 28, 684), 
(25, 23, 28, 26, 24, 22, 66, 72, 30, 21, 69, 29), 
(72, 30, 27, 69, 73, 31, 29, 25, 23, 74, 26, 66), 
(30, 32, 26, 28, 31, 33, 684, 679, 25, 35, 683, 27), 
(29, 28, 31, 32, 26, 27, 72, 74, 35, 25, 73, 33), 
(74, 35, 30, 73, 77, 36, 33, 29, 28, 80, 32, 72), 
(684, 29, 33, 686, 683, 26, 30, 35, 34, 679, 31, 687), 
(35, 34, 32, 31, 36, 37, 687, 684, 29, 38, 686, 30), 
(687, 33, 37, 691, 686, 32, 35, 38, 40, 684, 36, 692), 
(33, 31, 36, 34, 32, 30, 74, 80, 38, 29, 77, 37), 
(80, 38, 35, 77, 81, 39, 37, 33, 31, 82, 34, 74), 
(38, 40, 34, 36, 39, 41, 692, 687, 33, 43, 691, 35), 
(37, 36, 39, 40, 34, 35, 80, 82, 43, 33, 81, 41), 
(82, 43, 38, 81, 85, 44, 41, 37, 36, 88, 40, 80), 
(692, 37, 41, 694, 691, 34, 38, 43, 42, 687, 39, 695), 
(43, 42, 40, 39, 44, 45, 695, 692, 37, 46, 694, 38), 
(695, 41, 45, 699, 694, 40, 43, 46, 700, 692, 44, 700), 
(41, 39, 44, 42, 40, 38, 82, 88, 46, 37, 85, 45), 
(88, 46, 43, 85, 89, 47, 45, 41, 39, 90, 42, 82), 
(46, 700, 42, 44, 47, 702, 699, 695, 41, 703, 695, 43), 
(45, 44, 47, 700, 42, 43, 88, 90, 703, 41, 89, 702), 
(90, 703, 46, 89, 93, 707, 702, 45, 44, 708, 700, 88), 
(4, 152, 49, 6, 3, 149, 153, 51, 50, 146, 154, 7), 
(51, 50, 48, 154, 52, 53, 7, 4, 152, 54, 6, 153), 
(7, 49, 53, 11, 6, 48, 51, 54, 56, 4, 52, 12), 
(49, 154, 52, 50, 48, 153, 157, 96, 54, 152, 160, 53), 
(96, 54, 51, 160, 97, 55, 53, 49, 154, 98, 50, 157), 
(54, 56, 50, 52, 55, 57, 12, 7, 49, 59, 11, 51), 
(53, 52, 55, 56, 50, 51, 96, 98, 59, 49, 97, 57), 
(98, 59, 54, 97, 101, 60, 57, 53, 52, 104, 56, 96), 
(12, 53, 57, 14, 11, 50, 54, 59, 58, 7, 55, 15), 
(59, 58, 56, 55, 60, 61, 15, 12, 53, 62, 14, 54), 
(15, 57, 61, 19, 14, 56, 59, 62, 64, 12, 60, 20), 
(57, 55, 60, 58, 56, 54, 98, 104, 62, 53, 101, 61), 
(104, 62, 59, 101, 105, 63, 61, 57, 55, 106, 58, 98), 
(62, 64, 58, 60, 63, 65, 20, 15, 57, 67, 19, 59), 
(61, 60, 63, 64, 58, 59, 104, 106, 67, 57, 105, 65), 
(106, 67, 62, 105, 109, 68, 65, 61, 60, 112, 64, 104), 
(20, 61, 65, 22, 19, 58, 62, 67, 66, 15, 63, 23), 
(67, 66, 64, 63, 68, 69, 23, 20, 61, 70, 22, 62), 
(23, 65, 69, 27, 22, 64, 67, 70, 72, 20, 68, 28), 
(65, 63, 68, 66, 64, 62, 106, 112, 70, 61, 109, 69), 
(112, 70, 67, 109, 113, 71, 69, 65, 63, 114, 66, 106), 
(70, 72, 66, 68, 71, 73, 28, 23, 65, 75, 27, 67), 
(69, 68, 71, 72, 66, 67, 112, 114, 75, 65, 113, 73), 
(114, 75, 70, 113, 117, 76, 73, 69, 68, 120, 72, 112), 
(28, 69, 73, 30, 27, 66, 70, 75, 74, 23, 71, 31), 
(75, 74, 72, 71, 76, 77, 31, 28, 69, 78, 30, 70), 
(31, 73, 77, 35, 30, 72, 75, 78, 80, 28, 76, 36), 
(73, 71, 76, 74, 72, 70, 114, 120, 78, 69, 117, 77), 
(120, 78, 75, 117, 121, 79, 77, 73, 71, 122, 74, 114), 
(78, 80, 74, 76, 79, 81, 36, 31, 73, 83, 35, 75), 
(77, 76, 79, 80, 74, 75, 120, 122, 83, 73, 121, 81), 
(122, 83, 78, 121, 125, 84, 81, 77, 76, 128, 80, 120), 
(36, 77, 81, 38, 35, 74, 78, 83, 82, 31, 79, 39), 
(83, 82, 80, 79, 84, 85, 39, 36, 77, 86, 38, 78), 
(39, 81, 85, 43, 38, 80, 83, 86, 88, 36, 84, 44), 
(81, 79, 84, 82, 80, 78, 122, 128, 86, 77, 125, 85), 
(128, 86, 83, 125, 129, 87, 85, 81, 79, 130, 82, 122), 
(86, 88, 82, 84, 87, 89, 44, 39, 81, 91, 43, 83), 
(85, 84, 87, 88, 82, 83, 128, 130, 91, 81, 129, 89), 
(130, 91, 86, 129, 133, 92, 89, 85, 84, 136, 88, 128), 
(44, 85, 89, 46, 43, 82, 86, 91, 90, 39, 87, 47), 
(91, 90, 88, 87, 92, 93, 47, 44, 85, 94, 46, 86), 
(47, 89, 93, 703, 46, 88, 91, 94, 708, 44, 92, 707), 
(89, 87, 92, 90, 88, 86, 130, 136, 94, 85, 133, 93), 
(136, 94, 91, 133, 137, 95, 93, 89, 87, 138, 90, 130), 
(94, 708, 90, 92, 95, 710, 707, 47, 89, 711, 703, 91), 
(93, 92, 95, 708, 90, 91, 136, 138, 711, 89, 137, 710), 
(138, 711, 94, 137, 141, 715, 710, 93, 92, 716, 708, 136), 
(52, 160, 97, 54, 51, 157, 161, 99, 98, 154, 162, 55), 
(99, 98, 96, 162, 100, 101, 55, 52, 160, 102, 54, 161), 
(55, 97, 101, 59, 54, 96, 99, 102, 104, 52, 100, 60), 
(97, 162, 100, 98, 96, 161, 165, 168, 102, 160, 168, 101), 
(168, 102, 99, 165, 169, 103, 101, 97, 162, 170, 98, 162), 
(102, 104, 98, 100, 103, 105, 60, 55, 97, 107, 59, 99), 
(101, 100, 103, 104, 98, 99, 168, 170, 107, 97, 169, 105), 
(170, 107, 102, 169, 173, 108, 105, 101, 100, 176, 104, 168), 
(60, 101, 105, 62, 59, 98, 102, 107, 106, 55, 103, 63), 
(107, 106, 104, 103, 108, 109, 63, 60, 101, 110, 62, 102), 
(63, 105, 109, 67, 62, 104, 107, 110, 112, 60, 108, 68), 
(105, 103, 108, 106, 104, 102, 170, 176, 110, 101, 173, 109), 
(176, 110, 107, 173, 177, 111, 109, 105, 103, 178, 106, 170), 
(110, 112, 106, 108, 111, 113, 68, 63, 105, 115, 67, 107), 
(109, 108, 111, 112, 106, 107, 176, 178, 115, 105, 177, 113), 
(178, 115, 110, 177, 181, 116, 113, 109, 108, 184, 112, 176), 
(68, 109, 113, 70, 67, 106, 110, 115, 114, 63, 111, 71), 
(115, 114, 112, 111, 116, 117, 71, 68, 109, 118, 70, 110), 
(71, 113, 117, 75, 70, 112, 115, 118, 120, 68, 116, 76), 
(113, 111, 116, 114, 112, 110, 178, 184, 118, 109, 181, 117), 
(184, 118, 115, 181, 185, 119, 117, 113, 111, 186, 114, 178), 
(118, 120, 114, 116, 119, 121, 76, 71, 113, 123, 75, 115), 
(117, 116, 119, 120, 114, 115, 184, 186, 123, 113, 185, 121), 
(186, 123, 118, 185, 189, 124, 121, 117, 116, 124, 120, 184), 
(76, 117, 121, 78, 75, 114, 118, 123, 122, 71, 119, 79), 
(123, 122, 120, 119, 124, 125, 79, 76, 117, 126, 78, 118), 
(79, 121, 125, 83, 78, 120, 123, 126, 128, 76, 124, 84), 
(121, 119, 124, 122, 120, 118, 186, 189, 126, 117, 189, 125), 
(189, 126, 123, 186, 190, 127, 125, 121, 119, 191, 122, 119), 
(126, 128, 122, 124, 127, 129, 84, 79, 121, 131, 83, 123), 
(125, 124, 127, 128, 122, 123, 189, 191, 131, 121, 190, 129), 
(191, 131, 126, 190, 234, 132, 129, 125, 124, 237, 128, 189), 
(84, 125, 129, 86, 83, 122, 126, 131, 130, 79, 127, 87), 
(131, 130, 128, 127, 132, 133, 87, 84, 125, 134, 86, 126), 
(87, 129, 133, 91, 86, 128, 131, 134, 136, 84, 132, 92), 
(129, 127, 132, 130, 128, 126, 191, 237, 134, 125, 234, 133), 
(237, 134, 131, 234, 238, 135, 133, 129, 127, 239, 130, 191), 
(134, 136, 130, 132, 135, 137, 92, 87, 129, 139, 91, 131), 
(133, 132, 135, 136, 130, 131, 237, 239, 139, 129, 238, 137), 
(239, 139, 134, 238, 282, 140, 137, 133, 132, 285, 136, 237), 
(92, 133, 137, 94, 91, 130, 134, 139, 138, 87, 135, 95), 
(139, 138, 136, 135, 140, 141, 95, 92, 133, 142, 94, 134), 
(95, 137, 141, 711, 94, 136, 139, 142, 716, 92, 140, 715), 
(137, 135, 140, 138, 136, 134, 239, 285, 142, 133, 282, 141), 
(285, 142, 139, 282, 286, 143, 141, 137, 135, 287, 138, 239), 
(142, 716, 138, 140, 143, 718, 715, 95, 137, 719, 711, 139), 
(141, 140, 143, 716, 138, 139, 285, 287, 719, 137, 286, 718), 
(287, 719, 142, 286, 431, 575, 718, 141, 140, 287, 716, 285), 
(0, 288, 145, 1, 576, 432, 289, 147, 146, 0, 290, 3), 
(147, 146, 144, 290, 148, 149, 3, 0, 288, 150, 1, 289), 
(3, 145, 149, 4, 1, 144, 147, 150, 152, 0, 148, 48), 
(145, 290, 148, 146, 144, 289, 293, 192, 150, 288, 296, 149), 
(192, 150, 147, 296, 193, 151, 149, 145, 290, 194, 146, 293), 
(150, 152, 146, 148, 151, 153, 48, 3, 145, 155, 4, 147), 
(149, 148, 151, 152, 146, 147, 192, 194, 155, 145, 193, 153), 
(194, 155, 150, 193, 197, 156, 153, 149, 148, 200, 152, 192), 
(48, 149, 153, 49, 4, 146, 150, 155, 154, 3, 151, 51), 
(155, 154, 152, 151, 156, 157, 51, 48, 149, 158, 49, 150), 
(51, 153, 157, 52, 49, 152, 155, 158, 160, 48, 156, 96), 
(153, 151, 156, 154, 152, 150, 194, 200, 158, 149, 197, 157), 
(200, 158, 155, 197, 201, 159, 157, 153, 151, 202, 154, 194), 
(158, 160, 154, 156, 159, 161, 96, 51, 153, 163, 52, 155), 
(157, 156, 159, 160, 154, 155, 200, 202, 163, 153, 201, 161), 
(202, 163, 158, 201, 205, 164, 161, 157, 156, 208, 160, 200), 
(96, 157, 161, 97, 52, 154, 158, 163, 162, 51, 159, 99), 
(163, 162, 160, 159, 164, 165, 99, 96, 157, 166, 97, 158), 
(99, 161, 165, 100, 97, 160, 163, 166, 168, 96, 164, 168), 
(161, 159, 164, 162, 160, 158, 202, 208, 166, 157, 205, 165), 
(208, 166, 163, 205, 209, 167, 165, 161, 159, 210, 162, 202), 
(166, 168, 162, 164, 167, 169, 100, 99, 161, 171, 99, 163), 
(165, 164, 167, 168, 162, 163, 208, 210, 171, 161, 209, 169), 
(210, 171, 166, 209, 213, 172, 169, 165, 164, 216, 168, 208), 
(100, 165, 169, 102, 99, 162, 166, 171, 170, 162, 167, 103), 
(171, 170, 168, 167, 172, 173, 103, 100, 165, 174, 102, 166), 
(103, 169, 173, 107, 102, 168, 171, 174, 176, 100, 172, 108), 
(169, 167, 172, 170, 168, 166, 210, 216, 174, 165, 213, 173), 
(216, 174, 171, 213, 217, 175, 173, 169, 167, 218, 170, 210), 
(174, 176, 170, 172, 175, 177, 108, 103, 169, 179, 107, 171), 
(173, 172, 175, 176, 170, 171, 216, 218, 179, 169, 217, 177), 
(218, 179, 174, 217, 221, 180, 177, 173, 172, 224, 176, 216), 
(108, 173, 177, 110, 107, 170, 174, 179, 178, 103, 175, 111), 
(179, 178, 176, 175, 180, 181, 111, 108, 173, 182, 110, 174), 
(111, 177, 181, 115, 110, 176, 179, 182, 184, 108, 180, 116), 
(177, 175, 180, 178, 176, 174, 218, 224, 182, 173, 221, 181), 
(224, 182, 179, 221, 225, 183, 181, 177, 175, 226, 178, 218), 
(182, 184, 178, 180, 183, 185, 116, 111, 177, 187, 115, 179), 
(181, 180, 183, 184, 178, 179, 224, 226, 187, 177, 225, 185), 
(226, 187, 182, 225, 229, 188, 185, 181, 180, 232, 184, 224), 
(116, 181, 185, 118, 115, 178, 182, 187, 186, 111, 183, 119), 
(187, 186, 184, 183, 188, 189, 119, 116, 181, 190, 118, 182), 
(119, 185, 189, 123, 118, 184, 187, 190, 124, 116, 188, 124), 
(185, 183, 188, 186, 184, 182, 226, 232, 190, 181, 229, 189), 
(232, 190, 187, 229, 233, 191, 189, 185, 183, 234, 186, 226), 
(190, 124, 186, 188, 191, 126, 123, 119, 185, 127, 119, 187), 
(189, 188, 191, 124, 186, 187, 232, 234, 127, 185, 233, 126), 
(234, 127, 190, 233, 237, 131, 126, 189, 188, 132, 124, 232), 
(148, 296, 193, 150, 147, 293, 297, 195, 194, 290, 298, 151), 
(195, 194, 192, 298, 196, 197, 151, 148, 296, 198, 150, 297), 
(151, 193, 197, 155, 150, 192, 195, 198, 200, 148, 196, 156), 
(193, 298, 196, 194, 192, 297, 301, 240, 198, 296, 304, 197), 
(240, 198, 195, 304, 241, 199, 197, 193, 298, 242, 194, 301), 
(198, 200, 194, 196, 199, 201, 156, 151, 193, 203, 155, 195), 
(197, 196, 199, 200, 194, 195, 240, 242, 203, 193, 241, 201), 
(242, 203, 198, 241, 245, 204, 201, 197, 196, 248, 200, 240), 
(156, 197, 201, 158, 155, 194, 198, 203, 202, 151, 199, 159), 
(203, 202, 200, 199, 204, 205, 159, 156, 197, 206, 158, 198), 
(159, 201, 205, 163, 158, 200, 203, 206, 208, 156, 204, 164), 
(201, 199, 204, 202, 200, 198, 242, 248, 206, 197, 245, 205), 
(248, 206, 203, 245, 249, 207, 205, 201, 199, 250, 202, 242), 
(206, 208, 202, 204, 207, 209, 164, 159, 201, 211, 163, 203), 
(205, 204, 207, 208, 202, 203, 248, 250, 211, 201, 249, 209), 
(250, 211, 206, 249, 253, 212, 209, 205, 204, 256, 208, 248), 
(164, 205, 209, 166, 163, 202, 206, 211, 210, 159, 207, 167), 
(211, 210, 208, 207, 212, 213, 167, 164, 205, 214, 166, 206), 
(167, 209, 213, 171, 166, 208, 211, 214, 216, 164, 212, 172), 
(209, 207, 212, 210, 208, 206, 250, 256, 214, 205, 253, 213), 
(256, 214, 211, 253, 257, 215, 213, 209, 207, 258, 210, 250), 
(214, 216, 210, 212, 215, 217, 172, 167, 209, 219, 171, 211), 
(213, 212, 215, 216, 210, 211, 256, 258, 219, 209, 257, 217), 
(258, 219, 214, 257, 261, 220, 217, 213, 212, 264, 216, 256), 
(172, 213, 217, 174, 171, 210, 214, 219, 218, 167, 215, 175), 
(219, 218, 216, 215, 220, 221, 175, 172, 213, 222, 174, 214), 
(175, 217, 221, 179, 174, 216, 219, 222, 224, 172, 220, 180), 
(217, 215, 220, 218, 216, 214, 258, 264, 222, 213, 261, 221), 
(264, 222, 219, 261, 265, 223, 221, 217, 215, 266, 218, 258), 
(222, 224, 218, 220, 223, 225, 180, 175, 217, 227, 179, 219), 
(221, 220, 223, 224, 218, 219, 264, 266, 227, 217, 265, 225), 
(266, 227, 222, 265, 269, 228, 225, 221, 220, 272, 224, 264), 
(180, 221, 225, 182, 179, 218, 222, 227, 226, 175, 223, 183), 
(227, 226, 224, 223, 228, 229, 183, 180, 221, 230, 182, 222), 
(183, 225, 229, 187, 182, 224, 227, 230, 232, 180, 228, 188), 
(225, 223, 228, 226, 224, 222, 266, 272, 230, 221, 269, 229), 
(272, 230, 227, 269, 273, 231, 229, 225, 223, 274, 226, 266), 
(230, 232, 226, 228, 231, 233, 188, 183, 225, 235, 187, 227), 
(229, 228, 231, 232, 226, 227, 272, 274, 235, 225, 273, 233), 
(274, 235, 230, 273, 277, 236, 233, 229, 228, 280, 232, 272), 
(188, 229, 233, 190, 187, 226, 230, 235, 234, 183, 231, 191), 
(235, 234, 232, 231, 236, 237, 191, 188, 229, 238, 190, 230), 
(191, 233, 237, 127, 190, 232, 235, 238, 132, 188, 236, 131), 
(233, 231, 236, 234, 232, 230, 274, 280, 238, 229, 277, 237), 
(280, 238, 235, 277, 281, 239, 237, 233, 231, 282, 234, 274), 
(238, 132, 234, 236, 239, 134, 131, 191, 233, 135, 127, 235), 
(237, 236, 239, 132, 234, 235, 280, 282, 135, 233, 281, 134), 
(282, 135, 238, 281, 285, 139, 134, 237, 236, 140, 132, 280), 
(196, 304, 241, 198, 195, 301, 305, 243, 242, 298, 306, 199), 
(243, 242, 240, 306, 244, 245, 199, 196, 304, 246, 198, 305), 
(199, 241, 245, 203, 198, 240, 243, 246, 248, 196, 244, 204), 
(241, 306, 244, 242, 240, 305, 309, 312, 246, 304, 312, 245), 
(312, 246, 243, 309, 313, 247, 245, 241, 306, 314, 242, 306), 
(246, 248, 242, 244, 247, 249, 204, 199, 241, 251, 203, 243), 
(245, 244, 247, 248, 242, 243, 312, 314, 251, 241, 313, 249), 
(314, 251, 246, 313, 317, 252, 249, 245, 244, 320, 248, 312), 
(204, 245, 249, 206, 203, 242, 246, 251, 250, 199, 247, 207), 
(251, 250, 248, 247, 252, 253, 207, 204, 245, 254, 206, 246), 
(207, 249, 253, 211, 206, 248, 251, 254, 256, 204, 252, 212), 
(249, 247, 252, 250, 248, 246, 314, 320, 254, 245, 317, 253), 
(320, 254, 251, 317, 321, 255, 253, 249, 247, 322, 250, 314), 
(254, 256, 250, 252, 255, 257, 212, 207, 249, 259, 211, 251), 
(253, 252, 255, 256, 250, 251, 320, 322, 259, 249, 321, 257), 
(322, 259, 254, 321, 325, 260, 257, 253, 252, 328, 256, 320), 
(212, 253, 257, 214, 211, 250, 254, 259, 258, 207, 255, 215), 
(259, 258, 256, 255, 260, 261, 215, 212, 253, 262, 214, 254), 
(215, 257, 261, 219, 214, 256, 259, 262, 264, 212, 260, 220), 
(257, 255, 260, 258, 256, 254, 322, 328, 262, 253, 325, 261), 
(328, 262, 259, 325, 329, 263, 261, 257, 255, 330, 258, 322), 
(262, 264, 258, 260, 263, 265, 220, 215, 257, 267, 219, 259), 
(261, 260, 263, 264, 258, 259, 328, 330, 267, 257, 329, 265), 
(330, 267, 262, 329, 333, 268, 265, 261, 260, 268, 264, 328), 
(220, 261, 265, 222, 219, 258, 262, 267, 266, 215, 263, 223), 
(267, 266, 264, 263, 268, 269, 223, 220, 261, 270, 222, 262), 
(223, 265, 269, 227, 222, 264, 267, 270, 272, 220, 268, 228), 
(265, 263, 268, 266, 264, 262, 330, 333, 270, 261, 333, 269), 
(333, 270, 267, 330, 334, 271, 269, 265, 263, 335, 266, 263), 
(270, 272, 266, 268, 271, 273, 228, 223, 265, 275, 227, 267), 
(269, 268, 271, 272, 266, 267, 333, 335, 275, 265, 334, 273), 
(335, 275, 270, 334, 378, 276, 273, 269, 268, 381, 272, 333), 
(228, 269, 273, 230, 227, 266, 270, 275, 274, 223, 271, 231), 
(275, 274, 272, 271, 276, 277, 231, 228, 269, 278, 230, 270), 
(231, 273, 277, 235, 230, 272, 275, 278, 280, 228, 276, 236), 
(273, 271, 276, 274, 272, 270, 335, 381, 278, 269, 378, 277), 
(381, 278, 275, 378, 382, 279, 277, 273, 271, 383, 274, 335), 
(278, 280, 274, 276, 279, 281, 236, 231, 273, 283, 235, 275), 
(277, 276, 279, 280, 274, 275, 381, 383, 283, 273, 382, 281), 
(383, 283, 278, 382, 426, 284, 281, 277, 276, 429, 280, 381), 
(236, 277, 281, 238, 235, 274, 278, 283, 282, 231, 279, 239), 
(283, 282, 280, 279, 284, 285, 239, 236, 277, 286, 238, 278), 
(239, 281, 285, 135, 238, 280, 283, 286, 140, 236, 284, 139), 
(281, 279, 284, 282, 280, 278, 383, 429, 286, 277, 426, 285), 
(429, 286, 283, 426, 430, 287, 285, 281, 279, 431, 282, 383), 
(286, 140, 282, 284, 287, 142, 139, 239, 281, 143, 135, 283), 
(285, 284, 287, 140, 282, 283, 429, 431, 143, 281, 430, 142), 
(431, 143, 286, 430, 575, 719, 142, 285, 284, 431, 140, 429), 
(144, 432, 289, 145, 0, 576, 433, 291, 290, 144, 434, 147), 
(291, 290, 288, 434, 292, 293, 147, 144, 432, 294, 145, 433), 
(147, 289, 293, 148, 145, 288, 291, 294, 296, 144, 292, 192), 
(289, 434, 292, 290, 288, 433, 437, 336, 294, 432, 440, 293), 
(336, 294, 291, 440, 337, 295, 293, 289, 434, 338, 290, 437), 
(294, 296, 290, 292, 295, 297, 192, 147, 289, 299, 148, 291), 
(293, 292, 295, 296, 290, 291, 336, 338, 299, 289, 337, 297), 
(338, 299, 294, 337, 341, 300, 297, 293, 292, 344, 296, 336), 
(192, 293, 297, 193, 148, 290, 294, 299, 298, 147, 295, 195), 
(299, 298, 296, 295, 300, 301, 195, 192, 293, 302, 193, 294), 
(195, 297, 301, 196, 193, 296, 299, 302, 304, 192, 300, 240), 
(297, 295, 300, 298, 296, 294, 338, 344, 302, 293, 341, 301), 
(344, 302, 299, 341, 345, 303, 301, 297, 295, 346, 298, 338), 
(302, 304, 298, 300, 303, 305, 240, 195, 297, 307, 196, 299), 
(301, 300, 303, 304, 298, 299, 344, 346, 307, 297, 345, 305), 
(346, 307, 302, 345, 349, 308, 305, 301, 300, 352, 304, 344), 
(240, 301, 305, 241, 196, 298, 302, 307, 306, 195, 303, 243), 
(307, 306, 304, 303, 308, 309, 243, 240, 301, 310, 241, 302), 
(243, 305, 309, 244, 241, 304, 307, 310, 312, 240, 308, 312), 
(305, 303, 308, 306, 304, 302, 346, 352, 310, 301, 349, 309), 
(352, 310, 307, 349, 353, 311, 309, 305, 303, 354, 306, 346), 
(310, 312, 306, 308, 311, 313, 244, 243, 305, 315, 243, 307), 
(309, 308, 311, 312, 306, 307, 352, 354, 315, 305, 353, 313), 
(354, 315, 310, 353, 357, 316, 313, 309, 308, 360, 312, 352), 
(244, 309, 313, 246, 243, 306, 310, 315, 314, 306, 311, 247), 
(315, 314, 312, 311, 316, 317, 247, 244, 309, 318, 246, 310), 
(247, 313, 317, 251, 246, 312, 315, 318, 320, 244, 316, 252), 
(313, 311, 316, 314, 312, 310, 354, 360, 318, 309, 357, 317), 
(360, 318, 315, 357, 361, 319, 317, 313, 311, 362, 314, 354), 
(318, 320, 314, 316, 319, 321, 252, 247, 313, 323, 251, 315), 
(317, 316, 319, 320, 314, 315, 360, 362, 323, 313, 361, 321), 
(362, 323, 318, 361, 365, 324, 321, 317, 316, 368, 320, 360), 
(252, 317, 321, 254, 251, 314, 318, 323, 322, 247, 319, 255), 
(323, 322, 320, 319, 324, 325, 255, 252, 317, 326, 254, 318), 
(255, 321, 325, 259, 254, 320, 323, 326, 328, 252, 324, 260), 
(321, 319, 324, 322, 320, 318, 362, 368, 326, 317, 365, 325), 
(368, 326, 323, 365, 369, 327, 325, 321, 319, 370, 322, 362), 
(326, 328, 322, 324, 327, 329, 260, 255, 321, 331, 259, 323), 
(325, 324, 327, 328, 322, 323, 368, 370, 331, 321, 369, 329), 
(370, 331, 326, 369, 373, 332, 329, 325, 324, 376, 328, 368), 
(260, 325, 329, 262, 259, 322, 326, 331, 330, 255, 327, 263), 
(331, 330, 328, 327, 332, 333, 263, 260, 325, 334, 262, 326), 
(263, 329, 333, 267, 262, 328, 331, 334, 268, 260, 332, 268), 
(329, 327, 332, 330, 328, 326, 370, 376, 334, 325, 373, 333), 
(376, 334, 331, 373, 377, 335, 333, 329, 327, 378, 330, 370), 
(334, 268, 330, 332, 335, 270, 267, 263, 329, 271, 263, 331), 
(333, 332, 335, 268, 330, 331, 376, 378, 271, 329, 377, 270), 
(378, 271, 334, 377, 381, 275, 270, 333, 332, 276, 268, 376), 
(292, 440, 337, 294, 291, 437, 441, 339, 338, 434, 442, 295), 
(339, 338, 336, 442, 340, 341, 295, 292, 440, 342, 294, 441), 
(295, 337, 341, 299, 294, 336, 339, 342, 344, 292, 340, 300), 
(337, 442, 340, 338, 336, 441, 445, 384, 342, 440, 448, 341), 
(384, 342, 339, 448, 385, 343, 341, 337, 442, 386, 338, 445), 
(342, 344, 338, 340, 343, 345, 300, 295, 337, 347, 299, 339), 
(341, 340, 343, 344, 338, 339, 384, 386, 347, 337, 385, 345), 
(386, 347, 342, 385, 389, 348, 345, 341, 340, 392, 344, 384), 
(300, 341, 345, 302, 299, 338, 342, 347, 346, 295, 343, 303), 
(347, 346, 344, 343, 348, 349, 303, 300, 341, 350, 302, 342), 
(303, 345, 349, 307, 302, 344, 347, 350, 352, 300, 348, 308), 
(345, 343, 348, 346, 344, 342, 386, 392, 350, 341, 389, 349), 
(392, 350, 347, 389, 393, 351, 349, 345, 343, 394, 346, 386), 
(350, 352, 346, 348, 351, 353, 308, 303, 345, 355, 307, 347), 
(349, 348, 351, 352, 346, 347, 392, 394, 355, 345, 393, 353), 
(394, 355, 350, 393, 397, 356, 353, 349, 348, 400, 352, 392), 
(308, 349, 353, 310, 307, 346, 350, 355, 354, 303, 351, 311), 
(355, 354, 352, 351, 356, 357, 311, 308, 349, 358, 310, 350), 
(311, 353, 357, 315, 310, 352, 355, 358, 360, 308, 356, 316), 
(353, 351, 356, 354, 352, 350, 394, 400, 358, 349, 397, 357), 
(400, 358, 355, 397, 401, 359, 357, 353, 351, 402, 354, 394), 
(358, 360, 354, 356, 359, 361, 316, 311, 353, 363, 315, 355), 
(357, 356, 359, 360, 354, 355, 400, 402, 363, 353, 401, 361), 
(402, 363, 358, 401, 405, 364, 361, 357, 356, 408, 360, 400), 
(316, 357, 361, 318, 315, 354, 358, 363, 362, 311, 359, 319), 
(363, 362, 360, 359, 364, 365, 319, 316, 357, 366, 318, 358), 
(319, 361, 365, 323, 318, 360, 363, 366, 368, 316, 364, 324), 
(361, 359, 364, 362, 360, 358, 402, 408, 366, 357, 405, 365), 
(408, 366, 363, 405, 409, 367, 365, 361, 359, 410, 362, 402), 
(366, 368, 362, 364, 367, 369, 324, 319, 361, 371, 323, 363), 
(365, 364, 367, 368, 362, 363, 408, 410, 371, 361, 409, 369), 
(410, 371, 366, 409, 413, 372, 369, 365, 364, 416, 368, 408), 
(324, 365, 369, 326, 323, 362, 366, 371, 370, 319, 367, 327), 
(371, 370, 368, 367, 372, 373, 327, 324, 365, 374, 326, 366), 
(327, 369, 373, 331, 326, 368, 371, 374, 376, 324, 372, 332), 
(369, 367, 372, 370, 368, 366, 410, 416, 374, 365, 413, 373), 
(416, 374, 371, 413, 417, 375, 373, 369, 367, 418, 370, 410), 
(374, 376, 370, 372, 375, 377, 332, 327, 369, 379, 331, 371), 
(373, 372, 375, 376, 370, 371, 416, 418, 379, 369, 417, 377), 
(418, 379, 374, 417, 421, 380, 377, 373, 372, 424, 376, 416), 
(332, 373, 377, 334, 331, 370, 374, 379, 378, 327, 375, 335), 
(379, 378, 376, 375, 380, 381, 335, 332, 373, 382, 334, 374), 
(335, 377, 381, 271, 334, 376, 379, 382, 276, 332, 380, 275), 
(377, 375, 380, 378, 376, 374, 418, 424, 382, 373, 421, 381), 
(424, 382, 379, 421, 425, 383, 381, 377, 375, 426, 378, 418), 
(382, 276, 378, 380, 383, 278, 275, 335, 377, 279, 271, 379), 
(381, 380, 383, 276, 378, 379, 424, 426, 279, 377, 425, 278), 
(426, 279, 382, 425, 429, 283, 278, 381, 380, 284, 276, 424), 
(340, 448, 385, 342, 339, 445, 449, 387, 386, 442, 450, 343), 
(387, 386, 384, 450, 388, 389, 343, 340, 448, 390, 342, 449), 
(343, 385, 389, 347, 342, 384, 387, 390, 392, 340, 388, 348), 
(385, 450, 388, 386, 384, 449, 453, 456, 390, 448, 456, 389), 
(456, 390, 387, 453, 457, 391, 389, 385, 450, 458, 386, 450), 
(390, 392, 386, 388, 391, 393, 348, 343, 385, 395, 347, 387), 
(389, 388, 391, 392, 386, 387, 456, 458, 395, 385, 457, 393), 
(458, 395, 390, 457, 461, 396, 393, 389, 388, 464, 392, 456), 
(348, 389, 393, 350, 347, 386, 390, 395, 394, 343, 391, 351), 
(395, 394, 392, 391, 396, 397, 351, 348, 389, 398, 350, 390), 
(351, 393, 397, 355, 350, 392, 395, 398, 400, 348, 396, 356), 
(393, 391, 396, 394, 392, 390, 458, 464, 398, 389, 461, 397), 
(464, 398, 395, 461, 465, 399, 397, 393, 391, 466, 394, 458), 
(398, 400, 394, 396, 399, 401, 356, 351, 393, 403, 355, 395), 
(397, 396, 399, 400, 394, 395, 464, 466, 403, 393, 465, 401), 
(466, 403, 398, 465, 469, 404, 401, 397, 396, 472, 400, 464), 
(356, 397, 401, 358, 355, 394, 398, 403, 402, 351, 399, 359), 
(403, 402, 400, 399, 404, 405, 359, 356, 397, 406, 358, 398), 
(359, 401, 405, 363, 358, 400, 403, 406, 408, 356, 404, 364), 
(401, 399, 404, 402, 400, 398, 466, 472, 406, 397, 469, 405), 
(472, 406, 403, 469, 473, 407, 405, 401, 399, 474, 402, 466), 
(406, 408, 402, 404, 407, 409, 364, 359, 401, 411, 363, 403), 
(405, 404, 407, 408, 402, 403, 472, 474, 411, 401, 473, 409), 
(474, 411, 406, 473, 477, 412, 409, 405, 404, 412, 408, 472), 
(364, 405, 409, 366, 363, 402, 406, 411, 410, 359, 407, 367), 
(411, 410, 408, 407, 412, 413, 367, 364, 405, 414, 366, 406), 
(367, 409, 413, 371, 366, 408, 411, 414, 416, 364, 412, 372), 
(409, 407, 412, 410, 408, 406, 474, 477, 414, 405, 477, 413), 
(477, 414, 411, 474, 478, 415, 413, 409, 407, 479, 410, 407), 
(414, 416, 410, 412, 415, 417, 372, 367, 409, 419, 371, 411), 
(413, 412, 415, 416, 410, 411, 477, 479, 419, 409, 478, 417), 
(479, 419, 414, 478, 522, 420, 417, 413, 412, 525, 416, 477), 
(372, 413, 417, 374, 371, 410, 414, 419, 418, 367, 415, 375), 
(419, 418, 416, 415, 420, 421, 375, 372, 413, 422, 374, 414), 
(375, 417, 421, 379, 374, 416, 419, 422, 424, 372, 420, 380), 
(417, 415, 420, 418, 416, 414, 479, 525, 422, 413, 522, 421), 
(525, 422, 419, 522, 526, 423, 421, 417, 415, 527, 418, 479), 
(422, 424, 418, 420, 423, 425, 380, 375, 417, 427, 379, 419), 
(421, 420, 423, 424, 418, 419, 525, 527, 427, 417, 526, 425), 
(527, 427, 422, 526, 570, 428, 425, 421, 420, 573, 424, 525), 
(380, 421, 425, 382, 379, 418, 422, 427, 426, 375, 423, 383), 
(427, 426, 424, 423, 428, 429, 383, 380, 421, 430, 382, 422), 
(383, 425, 429, 279, 382, 424, 427, 430, 284, 380, 428, 283), 
(425, 423, 428, 426, 424, 422, 527, 573, 430, 421, 570, 429), 
(573, 430, 427, 570, 574, 431, 429, 425, 423, 575, 426, 527), 
(430, 284, 426, 428, 431, 286, 283, 383, 425, 287, 279, 427), 
(429, 428, 431, 284, 426, 427, 573, 575, 287, 425, 574, 286), 
(575, 287, 430, 574, 719, 143, 286, 429, 428, 575, 284, 573), 
(288, 576, 433, 289, 144, 0, 577, 435, 434, 288, 578, 291), 
(435, 434, 432, 578, 436, 437, 291, 288, 576, 438, 289, 577), 
(291, 433, 437, 292, 289, 432, 435, 438, 440, 288, 436, 336), 
(433, 578, 436, 434, 432, 577, 581, 480, 438, 576, 584, 437), 
(480, 438, 435, 584, 481, 439, 437, 433, 578, 482, 434, 581), 
(438, 440, 434, 436, 439, 441, 336, 291, 433, 443, 292, 435), 
(437, 436, 439, 440, 434, 435, 480, 482, 443, 433, 481, 441), 
(482, 443, 438, 481, 485, 444, 441, 437, 436, 488, 440, 480), 
(336, 437, 441, 337, 292, 434, 438, 443, 442, 291, 439, 339), 
(443, 442, 440, 439, 444, 445, 339, 336, 437, 446, 337, 438), 
(339, 441, 445, 340, 337, 440, 443, 446, 448, 336, 444, 384), 
(441, 439, 444, 442, 440, 438, 482, 488, 446, 437, 485, 445), 
(488, 446, 443, 485, 489, 447, 445, 441, 439, 490, 442, 482), 
(446, 448, 442, 444, 447, 449, 384, 339, 441, 451, 340, 443), 
(445, 444, 447, 448, 442, 443, 488, 490, 451, 441, 489, 449), 
(490, 451, 446, 489, 493, 452, 449, 445, 444, 496, 448, 488), 
(384, 445, 449, 385, 340, 442, 446, 451, 450, 339, 447, 387), 
(451, 450, 448, 447, 452, 453, 387, 384, 445, 454, 385, 446), 
(387, 449, 453, 388, 385, 448, 451, 454, 456, 384, 452, 456), 
(449, 447, 452, 450, 448, 446, 490, 496, 454, 445, 493, 453), 
(496, 454, 451, 493, 497, 455, 453, 449, 447, 498, 450, 490), 
(454, 456, 450, 452, 455, 457, 388, 387, 449, 459, 387, 451), 
(453, 452, 455, 456, 450, 451, 496, 498, 459, 449, 497, 457), 
(498, 459, 454, 497, 501, 460, 457, 453, 452, 504, 456, 496), 
(388, 453, 457, 390, 387, 450, 454, 459, 458, 450, 455, 391), 
(459, 458, 456, 455, 460, 461, 391, 388, 453, 462, 390, 454), 
(391, 457, 461, 395, 390, 456, 459, 462, 464, 388, 460, 396), 
(457, 455, 460, 458, 456, 454, 498, 504, 462, 453, 501, 461), 
(504, 462, 459, 501, 505, 463, 461, 457, 455, 506, 458, 498), 
(462, 464, 458, 460, 463, 465, 396, 391, 457, 467, 395, 459), 
(461, 460, 463, 464, 458, 459, 504, 506, 467, 457, 505, 465), 
(506, 467, 462, 505, 509, 468, 465, 461, 460, 512, 464, 504), 
(396, 461, 465, 398, 395, 458, 462, 467, 466, 391, 463, 399), 
(467, 466, 464, 463, 468, 469, 399, 396, 461, 470, 398, 462), 
(399, 465, 469, 403, 398, 464, 467, 470, 472, 396, 468, 404), 
(465, 463, 468, 466, 464, 462, 506, 512, 470, 461, 509, 469), 
(512, 470, 467, 509, 513, 471, 469, 465, 463, 514, 466, 506), 
(470, 472, 466, 468, 471, 473, 404, 399, 465, 475, 403, 467), 
(469, 468, 471, 472, 466, 467, 512, 514, 475, 465, 513, 473), 
(514, 475, 470, 513, 517, 476, 473, 469, 468, 520, 472, 512), 
(404, 469, 473, 406, 403, 466, 470, 475, 474, 399, 471, 407), 
(475, 474, 472, 471, 476, 477, 407, 404, 469, 478, 406, 470), 
(407, 473, 477, 411, 406, 472, 475, 478, 412, 404, 476, 412), 
(473, 471, 476, 474, 472, 470, 514, 520, 478, 469, 517, 477), 
(520, 478, 475, 517, 521, 479, 477, 473, 471, 522, 474, 514), 
(478, 412, 474, 476, 479, 414, 411, 407, 473, 415, 407, 475), 
(477, 476, 479, 412, 474, 475, 520, 522, 415, 473, 521, 414), 
(522, 415, 478, 521, 525, 419, 414, 477, 476, 420, 412, 520), 
(436, 584, 481, 438, 435, 581, 585, 483, 482, 578, 586, 439), 
(483, 482, 480, 586, 484, 485, 439, 436, 584, 486, 438, 585), 
(439, 481, 485, 443, 438, 480, 483, 486, 488, 436, 484, 444), 
(481, 586, 484, 482, 480, 585, 589, 528, 486, 584, 592, 485), 
(528, 486, 483, 592, 529, 487, 485, 481, 586, 530, 482, 589), 
(486, 488, 482, 484, 487, 489, 444, 439, 481, 491, 443, 483), 
(485, 484, 487, 488, 482, 483, 528, 530, 491, 481, 529, 489), 
(530, 491, 486, 529, 533, 492, 489, 485, 484, 536, 488, 528), 
(444, 485, 489, 446, 443, 482, 486, 491, 490, 439, 487, 447), 
(491, 490, 488, 487, 492, 493, 447, 444, 485, 494, 446, 486), 
(447, 489, 493, 451, 446, 488, 491, 494, 496, 444, 492, 452), 
(489, 487, 492, 490, 488, 486, 530, 536, 494, 485, 533, 493), 
(536, 494, 491, 533, 537, 495, 493, 489, 487, 538, 490, 530), 
(494, 496, 490, 492, 495, 497, 452, 447, 489, 499, 451, 491), 
(493, 492, 495, 496, 490, 491, 536, 538, 499, 489, 537, 497), 
(538, 499, 494, 537, 541, 500, 497, 493, 492, 544, 496, 536), 
(452, 493, 497, 454, 451, 490, 494, 499, 498, 447, 495, 455), 
(499, 498, 496, 495, 500, 501, 455, 452, 493, 502, 454, 494), 
(455, 497, 501, 459, 454, 496, 499, 502, 504, 452, 500, 460), 
(497, 495, 500, 498, 496, 494, 538, 544, 502, 493, 541, 501), 
(544, 502, 499, 541, 545, 503, 501, 497, 495, 546, 498, 538), 
(502, 504, 498, 500, 503, 505, 460, 455, 497, 507, 459, 499), 
(501, 500, 503, 504, 498, 499, 544, 546, 507, 497, 545, 505), 
(546, 507, 502, 545, 549, 508, 505, 501, 500, 552, 504, 544), 
(460, 501, 505, 462, 459, 498, 502, 507, 506, 455, 503, 463), 
(507, 506, 504, 503, 508, 509, 463, 460, 501, 510, 462, 502), 
(463, 505, 509, 467, 462, 504, 507, 510, 512, 460, 508, 468), 
(505, 503, 508, 506, 504, 502, 546, 552, 510, 501, 549, 509), 
(552, 510, 507, 549, 553, 511, 509, 505, 503, 554, 506, 546), 
(510, 512, 506, 508, 511, 513, 468, 463, 505, 515, 467, 507), 
(509, 508, 511, 512, 506, 507, 552, 554, 515, 505, 553, 513), 
(554, 515, 510, 553, 557, 516, 513, 509, 508, 560, 512, 552), 
(468, 509, 513, 470, 467, 506, 510, 515, 514, 463, 511, 471), 
(515, 514, 512, 511, 516, 517, 471, 468, 509, 518, 470, 510), 
(471, 513, 517, 475, 470, 512, 515, 518, 520, 468, 516, 476), 
(513, 511, 516, 514, 512, 510, 554, 560, 518, 509, 557, 517), 
(560, 518, 515, 557, 561, 519, 517, 513, 511, 562, 514, 554), 
(518, 520, 514, 516, 519, 521, 476, 471, 513, 523, 475, 515), 
(517, 516, 519, 520, 514, 515, 560, 562, 523, 513, 561, 521), 
(562, 523, 518, 561, 565, 524, 521, 517, 516, 568, 520, 560), 
(476, 517, 521, 478, 475, 514, 518, 523, 522, 471, 519, 479), 
(523, 522, 520, 519, 524, 525, 479, 476, 517, 526, 478, 518), 
(479, 521, 525, 415, 478, 520, 523, 526, 420, 476, 524, 419), 
(521, 519, 524, 522, 520, 518, 562, 568, 526, 517, 565, 525), 
(568, 526, 523, 565, 569, 527, 525, 521, 519, 570, 522, 562), 
(526, 420, 522, 524, 527, 422, 419, 479, 521, 423, 415, 523), 
(525, 524, 527, 420, 522, 523, 568, 570, 423, 521, 569, 422), 
(570, 423, 526, 569, 573, 427, 422, 525, 524, 428, 420, 568), 
(484, 592, 529, 486, 483, 589, 593, 531, 530, 586, 594, 487), 
(531, 530, 528, 594, 532, 533, 487, 484, 592, 534, 486, 593), 
(487, 529, 533, 491, 486, 528, 531, 534, 536, 484, 532, 492), 
(529, 594, 532, 530, 528, 593, 597, 600, 534, 592, 600, 533), 
(600, 534, 531, 597, 601, 535, 533, 529, 594, 602, 530, 594), 
(534, 536, 530, 532, 535, 537, 492, 487, 529, 539, 491, 531), 
(533, 532, 535, 536, 530, 531, 600, 602, 539, 529, 601, 537), 
(602, 539, 534, 601, 605, 540, 537, 533, 532, 608, 536, 600), 
(492, 533, 537, 494, 491, 530, 534, 539, 538, 487, 535, 495), 
(539, 538, 536, 535, 540, 541, 495, 492, 533, 542, 494, 534), 
(495, 537, 541, 499, 494, 536, 539, 542, 544, 492, 540, 500), 
(537, 535, 540, 538, 536, 534, 602, 608, 542, 533, 605, 541), 
(608, 542, 539, 605, 609, 543, 541, 537, 535, 610, 538, 602), 
(542, 544, 538, 540, 543, 545, 500, 495, 537, 547, 499, 539), 
(541, 540, 543, 544, 538, 539, 608, 610, 547, 537, 609, 545), 
(610, 547, 542, 609, 613, 548, 545, 541, 540, 616, 544, 608), 
(500, 541, 545, 502, 499, 538, 542, 547, 546, 495, 543, 503), 
(547, 546, 544, 543, 548, 549, 503, 500, 541, 550, 502, 542), 
(503, 545, 549, 507, 502, 544, 547, 550, 552, 500, 548, 508), 
(545, 543, 548, 546, 544, 542, 610, 616, 550, 541, 613, 549), 
(616, 550, 547, 613, 617, 551, 549, 545, 543, 618, 546, 610), 
(550, 552, 546, 548, 551, 553, 508, 503, 545, 555, 507, 547), 
(549, 548, 551, 552, 546, 547, 616, 618, 555, 545, 617, 553), 
(618, 555, 550, 617, 621, 556, 553, 549, 548, 556, 552, 616), 
(508, 549, 553, 510, 507, 546, 550, 555, 554, 503, 551, 511), 
(555, 554, 552, 551, 556, 557, 511, 508, 549, 558, 510, 550), 
(511, 553, 557, 515, 510, 552, 555, 558, 560, 508, 556, 516), 
(553, 551, 556, 554, 552, 550, 618, 621, 558, 549, 621, 557), 
(621, 558, 555, 618, 622, 559, 557, 553, 551, 623, 554, 551), 
(558, 560, 554, 556, 559, 561, 516, 511, 553, 563, 515, 555), 
(557, 556, 559, 560, 554, 555, 621, 623, 563, 553, 622, 561), 
(623, 563, 558, 622, 666, 564, 561, 557, 556, 669, 560, 621), 
(516, 557, 561, 518, 515, 554, 558, 563, 562, 511, 559, 519), 
(563, 562, 560, 559, 564, 565, 519, 516, 557, 566, 518, 558), 
(519, 561, 565, 523, 518, 560, 563, 566, 568, 516, 564, 524), 
(561, 559, 564, 562, 560, 558, 623, 669, 566, 557, 666, 565), 
(669, 566, 563, 666, 670, 567, 565, 561, 559, 671, 562, 623), 
(566, 568, 562, 564, 567, 569, 524, 519, 561, 571, 523, 563), 
(565, 564, 567, 568, 562, 563, 669, 671, 571, 561, 670, 569), 
(671, 571, 566, 670, 714, 572, 569, 565, 564, 717, 568, 669), 
(524, 565, 569, 526, 523, 562, 566, 571, 570, 519, 567, 527), 
(571, 570, 568, 567, 572, 573, 527, 524, 565, 574, 526, 566), 
(527, 569, 573, 423, 526, 568, 571, 574, 428, 524, 572, 427), 
(569, 567, 572, 570, 568, 566, 671, 717, 574, 565, 714, 573), 
(717, 574, 571, 714, 718, 575, 573, 569, 567, 719, 570, 671), 
(574, 428, 570, 572, 575, 430, 427, 527, 569, 431, 423, 571), 
(573, 572, 575, 428, 570, 571, 717, 719, 431, 569, 718, 430), 
(719, 431, 574, 718, 143, 287, 430, 573, 572, 719, 428, 717), 
(432, 0, 577, 433, 288, 144, 1, 579, 578, 432, 2, 435), 
(579, 578, 576, 2, 580, 581, 435, 432, 0, 582, 433, 1), 
(435, 577, 581, 436, 433, 576, 579, 582, 584, 432, 580, 480), 
(577, 2, 580, 578, 576, 1, 5, 624, 582, 0, 8, 581), 
(624, 582, 579, 8, 625, 583, 581, 577, 2, 626, 578, 5), 
(582, 584, 578, 580, 583, 585, 480, 435, 577, 587, 436, 579), 
(581, 580, 583, 584, 578, 579, 624, 626, 587, 577, 625, 585), 
(626, 587, 582, 625, 629, 588, 585, 581, 580, 632, 584, 624), 
(480, 581, 585, 481, 436, 578, 582, 587, 586, 435, 583, 483), 
(587, 586, 584, 583, 588, 589, 483, 480, 581, 590, 481, 582), 
(483, 585, 589, 484, 481, 584, 587, 590, 592, 480, 588, 528), 
(585, 583, 588, 586, 584, 582, 626, 632, 590, 581, 629, 589), 
(632, 590, 587, 629, 633, 591, 589, 585, 583, 634, 586, 626), 
(590, 592, 586, 588, 591, 593, 528, 483, 585, 595, 484, 587), 
(589, 588, 591, 592, 586, 587, 632, 634, 595, 585, 633, 593), 
(634, 595, 590, 633, 637, 596, 593, 589, 588, 640, 592, 632), 
(528, 589, 593, 529, 484, 586, 590, 595, 594, 483, 591, 531), 
(595, 594, 592, 591, 596, 597, 531, 528, 589, 598, 529, 590), 
(531, 593, 597, 532, 529, 592, 595, 598, 600, 528, 596, 600), 
(593, 591, 596, 594, 592, 590, 634, 640, 598, 589, 637, 597), 
(640, 598, 595, 637, 641, 599, 597, 593, 591, 642, 594, 634), 
(598, 600, 594, 596, 599, 601, 532, 531, 593, 603, 531, 595), 
(597, 596, 599, 600, 594, 595, 640, 642, 603, 593, 641, 601), 
(642, 603, 598, 641, 645, 604, 601, 597, 596, 648, 600, 640), 
(532, 597, 601, 534, 531, 594, 598, 603, 602, 594, 599, 535), 
(603, 602, 600, 599, 604, 605, 535, 532, 597, 606, 534, 598), 
(535, 601, 605, 539, 534, 600, 603, 606, 608, 532, 604, 540), 
(601, 599, 604, 602, 600, 598, 642, 648, 606, 597, 645, 605), 
(648, 606, 603, 645, 649, 607, 605, 601, 599, 650, 602, 642), 
(606, 608, 602, 604, 607, 609, 540, 535, 601, 611, 539, 603), 
(605, 604, 607, 608, 602, 603, 648, 650, 611, 601, 649, 609), 
(650, 611, 606, 649, 653, 612, 609, 605, 604, 656, 608, 648), 
(540, 605, 609, 542, 539, 602, 606, 611, 610, 535, 607, 543), 
(611, 610, 608, 607, 612, 613, 543, 540, 605, 614, 542, 606), 
(543, 609, 613, 547, 542, 608, 611, 614, 616, 540, 612, 548), 
(609, 607, 612, 610, 608, 606, 650, 656, 614, 605, 653, 613), 
(656, 614, 611, 653, 657, 615, 613, 609, 607, 658, 610, 650), 
(614, 616, 610, 612, 615, 617, 548, 543, 609, 619, 547, 611), 
(613, 612, 615, 616, 610, 611, 656, 658, 619, 609, 657, 617), 
(658, 619, 614, 657, 661, 620, 617, 613, 612, 664, 616, 656), 
(548, 613, 617, 550, 547, 610, 614, 619, 618, 543, 615, 551), 
(619, 618, 616, 615, 620, 621, 551, 548, 613, 622, 550, 614), 
(551, 617, 621, 555, 550, 616, 619, 622, 556, 548, 620, 556), 
(617, 615, 620, 618, 616, 614, 658, 664, 622, 613, 661, 621), 
(664, 622, 619, 661, 665, 623, 621, 617, 615, 666, 618, 658), 
(622, 556, 618, 620, 623, 558, 555, 551, 617, 559, 551, 619), 
(621, 620, 623, 556, 618, 619, 664, 666, 559, 617, 665, 558), 
(666, 559, 622, 665, 669, 563, 558, 621, 620, 564, 556, 664), 
(580, 8, 625, 582, 579, 5, 9, 627, 626, 2, 10, 583), 
(627, 626, 624, 10, 628, 629, 583, 580, 8, 630, 582, 9), 
(583, 625, 629, 587, 582, 624, 627, 630, 632, 580, 628, 588), 
(625, 10, 628, 626, 624, 9, 13, 672, 630, 8, 16, 629), 
(672, 630, 627, 16, 673, 631, 629, 625, 10, 674, 626, 13), 
(630, 632, 626, 628, 631, 633, 588, 583, 625, 635, 587, 627), 
(629, 628, 631, 632, 626, 627, 672, 674, 635, 625, 673, 633), 
(674, 635, 630, 673, 677, 636, 633, 629, 628, 680, 632, 672), 
(588, 629, 633, 590, 587, 626, 630, 635, 634, 583, 631, 591), 
(635, 634, 632, 631, 636, 637, 591, 588, 629, 638, 590, 630), 
(591, 633, 637, 595, 590, 632, 635, 638, 640, 588, 636, 596), 
(633, 631, 636, 634, 632, 630, 674, 680, 638, 629, 677, 637), 
(680, 638, 635, 677, 681, 639, 637, 633, 631, 682, 634, 674), 
(638, 640, 634, 636, 639, 641, 596, 591, 633, 643, 595, 635), 
(637, 636, 639, 640, 634, 635, 680, 682, 643, 633, 681, 641), 
(682, 643, 638, 681, 685, 644, 641, 637, 636, 688, 640, 680), 
(596, 637, 641, 598, 595, 634, 638, 643, 642, 591, 639, 599), 
(643, 642, 640, 639, 644, 645, 599, 596, 637, 646, 598, 638), 
(599, 641, 645, 603, 598, 640, 643, 646, 648, 596, 644, 604), 
(641, 639, 644, 642, 640, 638, 682, 688, 646, 637, 685, 645), 
(688, 646, 643, 685, 689, 647, 645, 641, 639, 690, 642, 682), 
(646, 648, 642, 644, 647, 649, 604, 599, 641, 651, 603, 643), 
(645, 644, 647, 648, 642, 643, 688, 690, 651, 641, 689, 649), 
(690, 651, 646, 689, 693, 652, 649, 645, 644, 696, 648, 688), 
(604, 645, 649, 606, 603, 642, 646, 651, 650, 599, 647, 607), 
(651, 650, 648, 647, 652, 653, 607, 604, 645, 654, 606, 646), 
(607, 649, 653, 611, 606, 648, 651, 654, 656, 604, 652, 612), 
(649, 647, 652, 650, 648, 646, 690, 696, 654, 645, 693, 653), 
(696, 654, 651, 693, 697, 655, 653, 649, 647, 698, 650, 690), 
(654, 656, 650, 652, 655, 657, 612, 607, 649, 659, 611, 651), 
(653, 652, 655, 656, 650, 651, 696, 698, 659, 649, 697, 657), 
(698, 659, 654, 697, 701, 660, 657, 653, 652, 704, 656, 696), 
(612, 653, 657, 614, 611, 650, 654, 659, 658, 607, 655, 615), 
(659, 658, 656, 655, 660, 661, 615, 612, 653, 662, 614, 654), 
(615, 657, 661, 619, 614, 656, 659, 662, 664, 612, 660, 620), 
(657, 655, 660, 658, 656, 654, 698, 704, 662, 653, 701, 661), 
(704, 662, 659, 701, 705, 663, 661, 657, 655, 706, 658, 698), 
(662, 664, 658, 660, 663, 665, 620, 615, 657, 667, 619, 659), 
(661, 660, 663, 664, 658, 659, 704, 706, 667, 657, 705, 665), 
(706, 667, 662, 705, 709, 668, 665, 661, 660, 712, 664, 704), 
(620, 661, 665, 622, 619, 658, 662, 667, 666, 615, 663, 623), 
(667, 666, 664, 663, 668, 669, 623, 620, 661, 670, 622, 662), 
(623, 665, 669, 559, 622, 664, 667, 670, 564, 620, 668, 563), 
(665, 663, 668, 666, 664, 662, 706, 712, 670, 661, 709, 669), 
(712, 670, 667, 709, 713, 671, 669, 665, 663, 714, 666, 706), 
(670, 564, 666, 668, 671, 566, 563, 623, 665, 567, 559, 667), 
(669, 668, 671, 564, 666, 667, 712, 714, 567, 665, 713, 566), 
(714, 567, 670, 713, 717, 571, 566, 669, 668, 572, 564, 712), 
(628, 16, 673, 630, 627, 13, 17, 675, 674, 10, 18, 631), 
(675, 674, 672, 18, 676, 677, 631, 628, 16, 678, 630, 17), 
(631, 673, 677, 635, 630, 672, 675, 678, 680, 628, 676, 636), 
(673, 18, 676, 674, 672, 17, 21, 24, 678, 16, 24, 677), 
(24, 678, 675, 21, 25, 679, 677, 673, 18, 26, 674, 18), 
(678, 680, 674, 676, 679, 681, 636, 631, 673, 683, 635, 675), 
(677, 676, 679, 680, 674, 675, 24, 26, 683, 673, 25, 681), 
(26, 683, 678, 25, 29, 684, 681, 677, 676, 32, 680, 24), 
(636, 677, 681, 638, 635, 674, 678, 683, 682, 631, 679, 639), 
(683, 682, 680, 679, 684, 685, 639, 636, 677, 686, 638, 678), 
(639, 681, 685, 643, 638, 680, 683, 686, 688, 636, 684, 644), 
(681, 679, 684, 682, 680, 678, 26, 32, 686, 677, 29, 685), 
(32, 686, 683, 29, 33, 687, 685, 681, 679, 34, 682, 26), 
(686, 688, 682, 684, 687, 689, 644, 639, 681, 691, 643, 683), 
(685, 684, 687, 688, 682, 683, 32, 34, 691, 681, 33, 689), 
(34, 691, 686, 33, 37, 692, 689, 685, 684, 40, 688, 32), 
(644, 685, 689, 646, 643, 682, 686, 691, 690, 639, 687, 647), 
(691, 690, 688, 687, 692, 693, 647, 644, 685, 694, 646, 686), 
(647, 689, 693, 651, 646, 688, 691, 694, 696, 644, 692, 652), 
(689, 687, 692, 690, 688, 686, 34, 40, 694, 685, 37, 693), 
(40, 694, 691, 37, 41, 695, 693, 689, 687, 42, 690, 34), 
(694, 696, 690, 692, 695, 697, 652, 647, 689, 699, 651, 691), 
(693, 692, 695, 696, 690, 691, 40, 42, 699, 689, 41, 697), 
(42, 699, 694, 41, 45, 700, 697, 693, 692, 700, 696, 40), 
(652, 693, 697, 654, 651, 690, 694, 699, 698, 647, 695, 655), 
(699, 698, 696, 695, 700, 701, 655, 652, 693, 702, 654, 694), 
(655, 697, 701, 659, 654, 696, 699, 702, 704, 652, 700, 660), 
(697, 695, 700, 698, 696, 694, 42, 45, 702, 693, 45, 701), 
(45, 702, 699, 42, 46, 703, 701, 697, 695, 47, 698, 695), 
(702, 704, 698, 700, 703, 705, 660, 655, 697, 707, 659, 699), 
(701, 700, 703, 704, 698, 699, 45, 47, 707, 697, 46, 705), 
(47, 707, 702, 46, 90, 708, 705, 701, 700, 93, 704, 45), 
(660, 701, 705, 662, 659, 698, 702, 707, 706, 655, 703, 663), 
(707, 706, 704, 703, 708, 709, 663, 660, 701, 710, 662, 702), 
(663, 705, 709, 667, 662, 704, 707, 710, 712, 660, 708, 668), 
(705, 703, 708, 706, 704, 702, 47, 93, 710, 701, 90, 709), 
(93, 710, 707, 90, 94, 711, 709, 705, 703, 95, 706, 47), 
(710, 712, 706, 708, 711, 713, 668, 663, 705, 715, 667, 707), 
(709, 708, 711, 712, 706, 707, 93, 95, 715, 705, 94, 713), 
(95, 715, 710, 94, 138, 716, 713, 709, 708, 141, 712, 93), 
(668, 709, 713, 670, 667, 706, 710, 715, 714, 663, 711, 671), 
(715, 714, 712, 711, 716, 717, 671, 668, 709, 718, 670, 710), 
(671, 713, 717, 567, 670, 712, 715, 718, 572, 668, 716, 571), 
(713, 711, 716, 714, 712, 710, 95, 141, 718, 709, 138, 717), 
(141, 718, 715, 138, 142, 719, 717, 713, 711, 143, 714, 95), 
(718, 572, 714, 716, 719, 574, 571, 671, 713, 575, 567, 715), 
(717, 716, 719, 572, 714, 715, 141, 143, 575, 713, 142, 574), 
(143, 575, 718, 142, 287, 431, 574, 717, 716, 143, 572, 141)	);


end Package_CB_Configuration;


package body Package_CB_Configuration is

end Package_CB_Configuration;